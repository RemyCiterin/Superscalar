import RvInstr::*;
import RvAlu::*;
import RvCSR::*;
