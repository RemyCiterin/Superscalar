import RvBranchPred :: *;
import Connectable :: *;
import BRAMCore :: *;
import RvICache :: *;
import TLTypes :: *;
import TLBram :: *;
import RvInstr :: *;
import Vector :: *;
import Assert :: *;
import Fifo :: *;

typedef struct {
  Super#(Bool) mask;
  Super#(Bit#(32)) uid;
  Super#(Bit#(32)) data;
  Super#(Bit#(32)) bprediction;
  Super#(CauseException) cause;
  Super#(Bool) exception;
  Super#(Bit#(32)) pc;
  Epoch epoch;
  BranchPredState bstate;
} FetchOutput deriving(Bits);

interface FetchIfc;
  method ActionValue#(FetchOutput) get;
  method Action redirect(Bit#(32) pc, Epoch newEpoch);

  method Action trainMis(BranchPredTrain infos);
  method Action trainHit(BranchPredTrain infos);

  interface TLMaster#(32, 32, 8, 8, 0) master;

  (* always_ready *) method Bit#(32) numMisPred;
endinterface

(* synthesize *)
module mkFetch(FetchIfc);
  Reg#(Epoch) nextEpoch[3] <- mkCReg(3, 0);
  Reg#(Bit#(32)) nextPc[3] <- mkCReg(3, 'h80000000);
  Reg#(Bit#(32)) uid <- mkReg(0);

  Bool bpredEnabled = True;

  ICache#(8, 8) icache <- mkICache(0);

  Fifo#(1, Tuple2#(Bit#(32), Epoch)) queue <- mkPipelineFifo;

  Bit#(32) pcMask = (1 << (supLogSize+2)) - 1;

  let bpred <- mkBranchPredictor;

  rule request;
    queue.enq(tuple2(nextPc[2], nextEpoch[2]));
    icache.lookup(nextPc[2] & ~pcMask);
    bpred.lookup(nextPc[2]);
  endrule

  interface master = icache.master;

  method numMisPred = bpred.numMisPred;

  method ActionValue#(FetchOutput) get if (queue.canDeq && icache.valid);
    match {.pc, .epoch} = queue.first;
    queue.deq;

    Bit#(32) currentUid = uid;
    Bit#(SupLogSize) laneBaseIndex = truncate(pc >> 2);
    Bit#(32) basePc = pc & ~pcMask;

    BranchPredState bstate = ?;
    Super#(Bool) mask = newVector;
    Super#(Bit#(32)) pcVec = newVector;
    Super#(Bit#(32)) uidVec = newVector;
    Super#(Bit#(32)) bprediction = newVector;
    for (Integer i=0; i < supSize; i = i + 1) begin
      Bool exception = False;
      mask[i] = exception ? fromInteger(i) == laneBaseIndex : fromInteger(i) >= laneBaseIndex;
      pcVec[i] = basePc + 4 * fromInteger(i);
      uidVec[i] = uid + fromInteger(i);
    end

    if (supLogSize == 0) mask[0] = True;

    if (epoch == nextEpoch[1]) begin
      match {.newPc, .offset, .bst} <- bpred.doPred();
      dynamicAssert(offset >= laneBaseIndex, "incoherent prediction");
      nextPc[1] <= bpredEnabled ? newPc : basePc + fromInteger(4*supSize);
      bstate = bst;

      for (Integer i=0; i < supSize; i = i + 1) begin
        bprediction[i] = supLogSize == 0 || offset == fromInteger(i) ? newPc : pcVec[i] + 4;
        if (bpredEnabled && offset < fromInteger(i) && supLogSize != 0) mask[i] = False;
        if (!bpredEnabled) bprediction[i] = pcVec[i] + 4;
      end
    end

    for (Integer i=0; i < supSize; i = i + 1) if (mask[i]) begin
      currentUid = currentUid + 1;
      uidVec[i] = currentUid;
    end

    icache.deq;

    uid <= currentUid;

    return FetchOutput {
      exception: replicate(False),
      cause: replicate(?),
      bprediction: bprediction,
      bstate: bstate,
      data: icache.response,
      epoch: epoch,
      uid: uidVec,
      mask: mask,
      pc: pcVec
    };
  endmethod

  method Action redirect(Bit#(32) newPc, Epoch newEpoch);
    nextEpoch[0] <= newEpoch;
    nextPc[0] <= newPc;
  endmethod

  method trainMis = bpred.trainMis;
  method trainHit = bpred.trainHit;
endmodule

typedef struct {
  Super#(Bool) mask;
  Super#(Bit#(32)) uid;
  Super#(RvInstr) instr;
  Super#(Bit#(32)) bprediction;
  Super#(CauseException) cause;
  BranchPredState bstate;
  Super#(Bool) exception;
  Super#(Bit#(32)) pc;
  Epoch epoch;
} Bundle deriving(Bits);

interface DecodeIfc;
  method Action put(FetchOutput in);
  method ActionValue#(Bundle) get;
  (* always_ready *) method Bool canGet;
endinterface

(* synthesize *)
module mkDecode(DecodeIfc);
  Fifo#(2, FetchOutput) fifo <- mkFifo;

  method Action put(FetchOutput in);
    fifo.enq(in);
  endmethod

  method canGet = fifo.canDeq;

  method ActionValue#(Bundle) get;
    let in = fifo.first;
    fifo.deq;

    Super#(RvInstr) instr = Vector::map(decodeRvInstr, in.data);
    Super#(CauseException) cause = in.cause;
    Super#(Bool) exception = in.exception;

    for (Integer i=0; i < supSize; i = i + 1) begin
      if (instr[i].opcode == Err && !exception[i]) begin
        cause[i] = IllegalInstruction;
        exception[i] = True;
      end
    end

    return Bundle{
      bprediction: in.bprediction,
      exception: exception,
      bstate: in.bstate,
      epoch: in.epoch,
      mask: in.mask,
      cause: cause,
      instr: instr,
      uid: in.uid,
      pc: in.pc
    };
  endmethod
endmodule

interface DispatchBuffer;
  // Give the current values inside the buffer
  (* always_ready *) method Bundle _read;

  // consume some values of the buffer, the values that we consumes mue be coherents:
  // if `0 <= a < b < supSize` are two indexes such that `self.mask[a] and self.mask[b]`, then we
  // can't consume `b` before consuming `a`, otherwise we may observe some data hazards...
  method Action consume(Super#(Bool) mask);

  // Read some values from the decode stage, only called if the fetch buffer is empty
  method Action put(Bundle in);
endinterface

module mkDispatchBuffer(DispatchBuffer);
  Reg#(Super#(Bool)) masks[2] <- mkCReg(2, replicate(False));
  Reg#(Super#(Bit#(32))) bpredictionBuf <- mkRegU;
  Reg#(Super#(CauseException)) causeBuf <- mkRegU;
  Reg#(Super#(Bool)) exceptionBuf <- mkRegU;
  Reg#(BranchPredState) bstateBuf <- mkRegU;
  Reg#(Super#(RvInstr)) instrBuf <- mkRegU;
  Reg#(Super#(Bit#(32))) uidBuf <- mkRegU;
  Reg#(Super#(Bit#(32))) pcBuf <- mkRegU;
  Reg#(Epoch) epochBuf <- mkRegU;

  method _read = Bundle{
    bprediction: bpredictionBuf,
    exception: exceptionBuf,
    bstate: bstateBuf,
    cause: causeBuf,
    instr: instrBuf,
    epoch: epochBuf,
    mask: masks[0],
    uid: uidBuf,
    pc: pcBuf
  };

  method Action consume(Super#(Bool) consumed);
    Super#(Bool) newMask = masks[0];
    Bool found = False;

    for (Integer i=0; i < supSize; i = i + 1) begin
      dynamicAssert(!found || !newMask[i] || !consumed[i], "DispatchBuffer<comsume> incoherent state");
      if (newMask[i] && !consumed[i]) found = True;
      if (consumed[i]) newMask[i] = False;
    end

    masks[0] <= newMask;
  endmethod

  method Action put(Bundle in) if (masks[1] == replicate(False));
    bpredictionBuf <= in.bprediction;
    exceptionBuf <= in.exception;
    bstateBuf <= in.bstate;
    instrBuf <= in.instr;
    epochBuf <= in.epoch;
    causeBuf <= in.cause;
    masks[1] <= in.mask;
    uidBuf <= in.uid;
    pcBuf <= in.pc;
  endmethod
endmodule

interface Buffer#(type t);
  // Give the current values inside the buffer
  (* always_ready *) method t _read;
  (* always_ready *) method Super#(Bool) mask;

  // consume some values of the buffer, the values that we consumes mue be coherents:
  // if `0 <= a < b < supSize` are two indexes such that `self.mask[a] and self.mask[b]`, then we
  // can't consume `b` before consuming `a`, otherwise we may observe some data hazards...
  method Action consume(Super#(Bool) msk);

  // Read some values from the decode stage, only called if the fetch buffer is empty
  method Action put(Super#(Bool) msk, t in);
endinterface

module mkBuffer(Buffer#(t)) provisos(Bits#(t, tW));
  Reg#(Super#(Bool)) masks[2] <- mkCReg(2, replicate(False));
  Reg#(t) value <- mkRegU;

  method _read = value;
  method mask = masks[0];

  method Action consume(Super#(Bool) consumed);
    Super#(Bool) newMask = masks[0];
    Bool found = False;

    for (Integer i=0; i < supSize; i = i + 1) begin
      dynamicAssert(!found || !newMask[i] || !consumed[i], "Buffer<comsume> incoherent state");
      if (newMask[i] && !consumed[i]) found = True;
      if (consumed[i]) newMask[i] = False;
    end

    masks[0] <= newMask;
  endmethod

  method Action put(Super#(Bool) msk, t in) if (masks[1] == replicate(False));
    masks[1] <= msk;
    value <= in;
  endmethod
endmodule
